module a (
    input logic  i_a
);

endmodule


module b (
    input logic  i_b
);

endmodule
//import td_pkg::* ;
import td_pkg::uvm_verbosity ;
import td_pkg::UVM_HIGH ;
module typedef_enum();

uvm_verbosity v;
initial begin
 v = UVM_HIGH;
end

endmodule


`define PRINT(STUFF) \
   begin \
       $display(STUFF);\
   end

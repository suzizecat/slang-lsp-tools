module a ();
typedef logic [10:2] my_type_t;
my_type_t  custom_type;

    logic a, b;

    assign a = b;


logic [31:0] an_array;

endmodule
import td_pkg::* ;
//import td_pkg::uvm_verbosity ;
module typedef_enum();

uvm_verbosity v;
initial begin
 v = UVM_HIGH;
end

endmodule

